`ifndef EVENT_UNIT_PKG
`define EVENT_UNIT_PKG


package event_unit_pkg;

    localparam logic        SIM                 = 1'b0;
    localparam logic        COVERGROUP_ANALYSIS = 1'b1;

endpackage


`endif
